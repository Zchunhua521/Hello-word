module
    initial begin
	    #1ns;
    end
endmodule
